module top_module(
    output zero
);

endmodule